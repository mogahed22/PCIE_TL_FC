module RX_main();
    buffer PD();
    buffer PH();
    buffer NPD();
    buffer NPH();
    buffer CD();
    buffer CH();
endmodule